  // I2C interface translator
